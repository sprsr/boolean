
// Module for Boolean Inverter Gate
// sprsr
////////////////////////////////////////////////
module INVERTER_GATE(input a, output y);
    assign y = !a;
endmodule
