// Module For Boolean XOR
//  @sprsr
////////////////////////////////////////////////////
module XOR_GATE(input a, input b, output y);
    assign y = a ^ b; 
endmodule
