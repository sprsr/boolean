# Module for Boolean AND Gate
# sprsr
#######################################################
module AND_GATE(input a, input b, output y);
    assign y = a & b;
end module
